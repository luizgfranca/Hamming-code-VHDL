LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HAMMING_SENDER IS
	PORT (ENTRADA : IN STD_LOGIC_VECTOR(8 DOWNTO 1);
			SAIDA : OUT STD_LOGIC_VECTOR(12 DOWNTO 1) );
END HAMMING_SENDER;

ARCHITECTURE SENDER OF HAMMING_SENDER IS
BEGIN	
	-- PRIMEIRAMENTE COLOCO OS BITS DA MENSAGEM NA POSIÇÃO CERTA
	SAIDA(3) <= ENTRADA(1);
	SAIDA(5) <= ENTRADA(2);
	SAIDA(6) <= ENTRADA(3);
	SAIDA(7) <= ENTRADA(4);
	SAIDA(9) <= ENTRADA(5);
	SAIDA(10) <= ENTRADA(6);
	SAIDA(11) <= ENTRADA(7);
	SAIDA(12) <= ENTRADA(8);
	
	-- AGORA CALCULO OS BITS DE PARIDADE
	SAIDA(1) <= ENTRADA(1) XOR ENTRADA(2) XOR ENTRADA(4) XOR ENTRADA(5) XOR ENTRADA(7);
	SAIDA(2) <= ENTRADA(1) XOR ENTRADA(3) XOR ENTRADA(4) XOR ENTRADA(6) XOR ENTRADA(7);
	SAIDA(4) <= ENTRADA(2) XOR ENTRADA(3) XOR ENTRADA(4) XOR ENTRADA(8);
	SAIDA(8) <= ENTRADA(5) XOR ENTRADA(6) XOR ENTRADA(7) XOR ENTRADA(8);

END SENDER;